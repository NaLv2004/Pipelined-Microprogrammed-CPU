 module CPUTop0000000001 ;
 reg clk;
 reg rst;
 wire [15:0] imem_addr;
 wire [31:0] imem_data;
 wire [7:0] register_file_addr_1;
 wire [7:0] register_file_addr_2;
 wire [15:0] register_data_out_1;
 wire [15:0] register_data_out_2;
 wire [31:0] micro_code;
 wire [7:0] micro_code_addr;
 wire [31:0] micro_code_speculative_fetch;  // REASSIGN!
 wire [7:0] micro_code_addr_speculative_fetch;  // REASSIGN!
 wire [15:0] alu_result;
 wire [15:0] data_memory_alu;
 wire [7:0] address_memory_alu;
 wire [0:0] write_en_memory;
 wire [0:0] write_en_regfile;
 wire [7:0] register_file_addr_dest;
 wire [15:0] mem_regfile_test;
 wire [15:0] mem_external_test;
 wire [15:0] mem_regfile_test1;
 wire [15:0] mem_external_test1;
 wire [0:0] flush_pipeline; // flush pipeline when branch prediction fails
 wire dec_ready;
 wire exec_ready; // connects CU and Fetch
 // fe-de; de-cu; cu-alu; alu-fe interfaces
 wire [49:0] fetch_idecode_interface;
 wire [91:0] idecode_cu_interface;
 wire [112:0] cu_alu_interface;
 wire [18:0] alu_fetch_interface;
 wire [31:0] micro_code_cu_external_mem;
 assign mem_regfile_test1 = u_0000000001_RegisterFile0000000001.mem[1];
 assign mem_external_test1 = u_0000000001_ExternalMem0000000001.mem[1];
Fetch0000000001  u_0000000001_Fetch0000000001(.clk(clk), .rst(rst), .imem_addr(imem_addr), .imem_data(imem_data), .dec_ready(dec_ready), .exec_ready(exec_ready), .flush_pipeline(flush_pipeline), .fetch_idecode_interface(fetch_idecode_interface), .alu_fetch_interface(alu_fetch_interface));
InstrMem0000000001  u_0000000001_InstrMem0000000001(.addr(imem_addr), .data_out(imem_data));
Decode0000000001  u_0000000001_Decode0000000001(.clk(clk), .rst(rst), .dec_ready(dec_ready), .flush_pipeline(flush_pipeline), .fetch_idecode_interface(fetch_idecode_interface), .idecode_cu_interface(idecode_cu_interface));
CU0000000001  u_0000000001_CU0000000001(.clk(clk), .rst(rst), .micro_code_in_normal(micro_code), .micro_code_in_speculative(micro_code_speculative_fetch), .micro_code_addr_out(micro_code_addr), .micro_code_addr_speculative_fetch(micro_code_addr_speculative_fetch), .o_exec_ready_combined(exec_ready), .flush_pipeline(flush_pipeline), .idecode_cu_interface(idecode_cu_interface), .cu_alu_interface(cu_alu_interface), .micro_code_out_external_mem(micro_code_cu_external_mem));
RegisterFile0000000001  u_0000000001_RegisterFile0000000001(.clk(clk), .reg_addr_1(register_file_addr_1), .reg_addr_2(register_file_addr_2), .data_out_1(register_data_out_1), .data_out_2(register_data_out_2), .write_en(write_en_regfile), .reg_addr_in(register_file_addr_dest), .data_in(alu_result), .mem_test(mem_regfile_test));
MicroInstrMem0000000001  u_0000000001_MicroInstrMem0000000001(.micro_code_addr_in(micro_code_addr), .micro_code_data_out(micro_code), .micro_code_addr_speculative_fetch_in(micro_code_addr_speculative_fetch), .micro_code_data_speculative_fetch_out(micro_code_speculative_fetch));
ExternalMem0000000001  u_0000000001_ExternalMem0000000001(.clk(clk), .micro_code(micro_code_cu_external_mem), .addr(address_memory_alu), .data_in(alu_result), .data_out(data_memory_alu), .data_test(mem_external_test));
ALU0000000001  u_0000000001_ALU0000000001(.clk(clk), .alu_regfile_in_1(register_data_out_1), .alu_regfile_in_2(register_data_out_2), .alu_memory_in(data_memory_alu), .alu_result(alu_result), .alu_regfile_address_out_1(register_file_addr_1), .alu_regfile_address_out_2(register_file_addr_2), .alu_memory_address_out(address_memory_alu), .alu_memory_write_en_out(write_en_memory), .alu_regfile_write_en_out(write_en_regfile), .alu_regfile_address_out(register_file_addr_dest), .cu_alu_interface(cu_alu_interface), .alu_fetch_interface(alu_fetch_interface));
 always #5 clk = ~clk;
 initial begin
   clk = 0;
   rst = 1;
   #10 rst = 0;
 end
 initial begin
 u_0000000001_InstrMem0000000001.mem[0] = 32'b10000000_00001000_00000000_00000000;
 u_0000000001_InstrMem0000000001.mem[1] = 32'b10000000_00000101_00000000_00000001;
 u_0000000001_InstrMem0000000001.mem[2] = 32'b00000001_00000001_00000010_00000000;
 u_0000000001_InstrMem0000000001.mem[3] = 32'b00100001_00000001_00001010_00000000;
 u_0000000001_InstrMem0000000001.mem[4] = 32'b10000001_00000000_00000000_00000000;
 u_0000000001_InstrMem0000000001.mem[5] = 32'b00010001_00000001_00000011_00000001;
 u_0000000001_InstrMem0000000001.mem[6] = 32'b00100010_00000001_00000001_00000001;
 u_0000000001_InstrMem0000000001.mem[7] = 32'b00100001_00000001_00001010_00000001;
 u_0000000001_InstrMem0000000001.mem[8] = 32'b10000000_00000001_00000000_00000100;
 u_0000000001_InstrMem0000000001.mem[9] = 32'b10000001_00000001_00000001_00000000;
 u_0000000001_InstrMem0000000001.mem[10] = 32'b00100001_00000000_00010000_00000000;
 u_0000000001_InstrMem0000000001.mem[11] = 32'b01100000_00000000_00000001_00001000;
 u_0000000001_InstrMem0000000001.mem[12] = 32'b10000001_00000001_00000010_00000000;
 // ['add rd, rs1, rs2'];
 u_0000000001_MicroInstrMem0000000001.mem[0] = 16'b0001000011000001;
 // ['sub rd, rs1, rs2'];
 u_0000000001_MicroInstrMem0000000001.mem[1] = 16'b0010000011000001;
 // ['and rd, rs1, rs2'];
 u_0000000001_MicroInstrMem0000000001.mem[2] = 16'b0011000011000001;
 // ['or rd, rs1, rs2'];
 u_0000000001_MicroInstrMem0000000001.mem[3] = 16'b0100000011000001;
 // ['xor rd, rs1, rs2'];
 u_0000000001_MicroInstrMem0000000001.mem[4] = 16'b0101000011000001;
 // ['sll rd, rs1, rs2'];
 u_0000000001_MicroInstrMem0000000001.mem[5] = 16'b0110000011000001;
 // ['srl rd, rs1, rs2'];
 u_0000000001_MicroInstrMem0000000001.mem[6] = 16'b0111000011000001;
 // ['add rd, [mem1], rs2'];
 u_0000000001_MicroInstrMem0000000001.mem[7] = 20'b00100000100000010000;
 u_0000000001_MicroInstrMem0000000001.mem[8] = 20'b00000000000000001000;
 u_0000000001_MicroInstrMem0000000001.mem[9] = 20'b00010001001001000001;
 // ['add rd, rs1, [mem2]'];
 u_0000000001_MicroInstrMem0000000001.mem[10] = 20'b00100000010000010000;
 u_0000000001_MicroInstrMem0000000001.mem[11] = 20'b00000000000000001000;
 u_0000000001_MicroInstrMem0000000001.mem[12] = 20'b00010001000110000001;
 // ['sub rd, [mem1], rs2'];
 u_0000000001_MicroInstrMem0000000001.mem[13] = 20'b00100000100000010000;
 u_0000000001_MicroInstrMem0000000001.mem[14] = 20'b00000000000000001000;
 u_0000000001_MicroInstrMem0000000001.mem[15] = 20'b00010010001001000001;
 // ['sub rd, rs1, [mem2]'];
 u_0000000001_MicroInstrMem0000000001.mem[16] = 20'b00100000010000010000;
 u_0000000001_MicroInstrMem0000000001.mem[17] = 20'b00000000000000001000;
 u_0000000001_MicroInstrMem0000000001.mem[18] = 20'b00010010000110000001;
 // ['and rd, [mem1], rs2'];
 u_0000000001_MicroInstrMem0000000001.mem[19] = 20'b00100000100000010000;
 u_0000000001_MicroInstrMem0000000001.mem[20] = 20'b00000000000000001000;
 u_0000000001_MicroInstrMem0000000001.mem[21] = 20'b00010011001001000001;
 // ['and rd, rs1, [mem2]'];
 u_0000000001_MicroInstrMem0000000001.mem[22] = 20'b00100000010000010000;
 u_0000000001_MicroInstrMem0000000001.mem[23] = 20'b00000000000000001000;
 u_0000000001_MicroInstrMem0000000001.mem[24] = 20'b00010011000110000001;
 // ['or rd, [mem1], rs2'];
 u_0000000001_MicroInstrMem0000000001.mem[25] = 20'b00100000100000010000;
 u_0000000001_MicroInstrMem0000000001.mem[26] = 20'b00000000000000001000;
 u_0000000001_MicroInstrMem0000000001.mem[27] = 20'b00010100001001000001;
 // ['or rd, rs1, [mem2]'];
 u_0000000001_MicroInstrMem0000000001.mem[28] = 20'b00100000010000010000;
 u_0000000001_MicroInstrMem0000000001.mem[29] = 20'b00000000000000001000;
 u_0000000001_MicroInstrMem0000000001.mem[30] = 20'b00010100000110000001;
 // ['xor rd, [mem1], rs2'];
 u_0000000001_MicroInstrMem0000000001.mem[31] = 20'b00100000100000010000;
 u_0000000001_MicroInstrMem0000000001.mem[32] = 20'b00000000000000001000;
 u_0000000001_MicroInstrMem0000000001.mem[33] = 20'b00010101001001000001;
 // ['xor rd, rs1, [mem2]'];
 u_0000000001_MicroInstrMem0000000001.mem[34] = 20'b00100000010000010000;
 u_0000000001_MicroInstrMem0000000001.mem[35] = 20'b00000000000000001000;
 u_0000000001_MicroInstrMem0000000001.mem[36] = 20'b00010101000110000001;
 // ['sll rd, [mem1], rs2'];
 u_0000000001_MicroInstrMem0000000001.mem[37] = 20'b00100000100000010000;
 u_0000000001_MicroInstrMem0000000001.mem[38] = 20'b00000000000000001000;
 u_0000000001_MicroInstrMem0000000001.mem[39] = 20'b00010110001001000001;
 // ['sll rd, rs1, [mem2]'];
 u_0000000001_MicroInstrMem0000000001.mem[40] = 20'b00100000010000010000;
 u_0000000001_MicroInstrMem0000000001.mem[41] = 20'b00000000000000001000;
 u_0000000001_MicroInstrMem0000000001.mem[42] = 20'b00010110000110000001;
 // ['srl rd, [mem1], rs2'];
 u_0000000001_MicroInstrMem0000000001.mem[43] = 20'b00100000100000010000;
 u_0000000001_MicroInstrMem0000000001.mem[44] = 20'b00000000000000001000;
 u_0000000001_MicroInstrMem0000000001.mem[45] = 20'b00010111001001000001;
 // ['srl rd, rs1, [mem2]'];
 u_0000000001_MicroInstrMem0000000001.mem[46] = 20'b00100000010000010000;
 u_0000000001_MicroInstrMem0000000001.mem[47] = 20'b00000000000000001000;
 u_0000000001_MicroInstrMem0000000001.mem[48] = 20'b00010111000110000001;
 // ['add rd, rs1, imm'];
 u_0000000001_MicroInstrMem0000000001.mem[49] = 21'b100000001000010000001;
 // ['sub rd, rs1, imm'];
 u_0000000001_MicroInstrMem0000000001.mem[50] = 21'b100000010000010000001;
 // ['and rd, rs1, imm'];
 u_0000000001_MicroInstrMem0000000001.mem[51] = 21'b100000011000010000001;
 // ['or rd, rs1, imm'];
 u_0000000001_MicroInstrMem0000000001.mem[52] = 21'b100000100000010000001;
 // ['xor rd, rs1, imm'];
 u_0000000001_MicroInstrMem0000000001.mem[53] = 21'b100000101000010000001;
 // ['sll rd, rs1, imm'];
 u_0000000001_MicroInstrMem0000000001.mem[54] = 21'b100000110000010000001;
 // ['srl rd, rs1, imm'];
 u_0000000001_MicroInstrMem0000000001.mem[55] = 21'b100000111000010000001;
 // ['jump imm'];
 u_0000000001_MicroInstrMem0000000001.mem[56] = 16'b0000000000000000;
 // ['beq rs1, rs2, imm'];
 u_0000000001_MicroInstrMem0000000001.mem[57] = 16'b1100000011000000;
 // ['load rd, [mem1]'];
 u_0000000001_MicroInstrMem0000000001.mem[58] = 20'b00100000100000010000;
 u_0000000001_MicroInstrMem0000000001.mem[59] = 20'b000000001000;
 u_0000000001_MicroInstrMem0000000001.mem[60] = 20'b00010000001000000001;
 // ['store [mem1], rs1'];
 u_0000000001_MicroInstrMem0000000001.mem[61] = 16'b0000_0100_1001_0100;
 u_0000000001_MicroInstrMem0000000001.mem[62] = 16'b0000_0000_0000_0010;
 // ['store [mem1], imm'];
 u_0000000001_MicroInstrMem0000000001.mem[63] = 22'b10_0000_0000_0100_0001_0100;
 u_0000000001_MicroInstrMem0000000001.mem[64] = 16'b0000_0000_0000_0010;
 // ['NO-OP(Used when flushing pipeline)'];
 u_0000000001_MicroInstrMem0000000001.mem[65] = 16'b0000000000000000;
 u_0000000001_MicroInstrMem0000000001.mem[255] = 16'b0000_0000;
 u_0000000001_ExternalMem0000000001.mem[0] = 16'b0000_0001;
 u_0000000001_ExternalMem0000000001.mem[1] = 16'b0001_0010;
 u_0000000001_ExternalMem0000000001.mem[2] = 16'b0010_0000;
 u_0000000001_ExternalMem0000000001.mem[3] = 16'b0000_0100;
 u_0000000001_ExternalMem0000000001.mem[4] = 16'b0000_0101;
 u_0000000001_ExternalMem0000000001.mem[5] = 16'b0000_0110;
 u_0000000001_ExternalMem0000000001.mem[6] = 16'b0000_0111;
 u_0000000001_ExternalMem0000000001.mem[7] = 16'b0000_1000;
 u_0000000001_ExternalMem0000000001.mem[8] = 16'b0000_1111;
 u_0000000001_ExternalMem0000000001.mem[9] = 16'b0000_1010;
 u_0000000001_ExternalMem0000000001.mem[10] = 16'b0000_1011;
 u_0000000001_RegisterFile0000000001.mem[0] = 16'b0000_0000_0000_0001;
 u_0000000001_RegisterFile0000000001.mem[1] = 16'b0000_0000_0000_0010;
 u_0000000001_RegisterFile0000000001.mem[2] = 16'b0000_0000_0000_0011;
 u_0000000001_RegisterFile0000000001.mem[3] = 16'b0000_0000_0000_0101;
 u_0000000001_RegisterFile0000000001.mem[4] = 16'b0000_0000_0000_0110;
 u_0000000001_RegisterFile0000000001.mem[5] = 16'b0000_0000_0000_0111;
 u_0000000001_RegisterFile0000000001.mem[6] = 16'b0000_0000_0000_1000;
 u_0000000001_RegisterFile0000000001.mem[7] = 16'b0000_0000_0000_1001;
 u_0000000001_RegisterFile0000000001.mem[8] = 16'b0000_0000_0000_1010;
 u_0000000001_RegisterFile0000000001.mem[9] = 16'b0000_0000_0000_1011;
 u_0000000001_RegisterFile0000000001.mem[10] = 16'b0000_0000_0000_1100;
 u_0000000001_RegisterFile0000000001.mem[11] = 16'b0000_0000_0000_1101;
 u_0000000001_RegisterFile0000000001.mem[12] = 16'b0000_0000_0000_1110;
 u_0000000001_RegisterFile0000000001.mem[13] = 16'b0000_0000_0000_1111;
 u_0000000001_RegisterFile0000000001.mem[14] = 16'b0000_0000_0001_0000;
 u_0000000001_RegisterFile0000000001.mem[15] = 16'b0000_0000_0001_0001;
 u_0000000001_RegisterFile0000000001.mem[16] = 16'b0000_0000_0001_0010;
 u_0000000001_RegisterFile0000000001.mem[17] = 16'b0000_0000_0001_0011;
 end
 initial begin
     $dumpfile("wave.vcd");
     $dumpvars(0, CPUTop0000000001);
     #2500
     $finish;
 end
 endmodule
